// ================================================================
// NVDLA Open Source Project
//
// Copyright(c) 2016 - 2017 NVIDIA Corporation. Licensed under the
// NVDLA Open Hardware License; Check "LICENSE" which comes with
// this distribution for more information.
// ================================================================
// File Name: NV_NVDLA_SDP_HLS_X_int_mul.v
module NV_NVDLA_SDP_HLS_X_int_mul (
   alu_data_out //|< i
  ,alu_out_pvld //|< i
  ,cfg_mul_bypass //|< i
  ,cfg_mul_op //|< i
  ,cfg_mul_prelu //|< i
  ,cfg_mul_src //|< i
  ,chn_mul_op //|< i
  ,mul_op_pvld //|< i
  ,mul_out_prdy //|< i
  ,nvdla_core_clk //|< i
  ,nvdla_core_rstn //|< i
  ,alu_out_prdy //|> o
  ,bypass_trt_out //|> o
  ,mul_data_out //|> o
  ,mul_op_prdy //|> o
  ,mul_out_pvld //|> o
  );
input [32:0] alu_data_out;
input alu_out_pvld;
input cfg_mul_bypass;
input [15:0] cfg_mul_op;
input cfg_mul_prelu;
input cfg_mul_src;
input [15:0] chn_mul_op;
input mul_op_pvld;
input mul_out_prdy;
input nvdla_core_clk;
input nvdla_core_rstn;
output alu_out_prdy;
output bypass_trt_out;
output [48:0] mul_data_out;
output mul_op_prdy;
output mul_out_pvld;
wire alu_out_srdy;
wire bypass_trt;
wire bypass_trt_reg;
wire [48:0] mul_data_final;
wire [32:0] mul_data_in;
wire [32:0] mul_data_sync;
wire mul_final_prdy;
wire mul_final_pvld;
wire [15:0] mul_op_in;
wire [15:0] mul_op_sync;
wire [48:0] mul_prelu_out;
wire mul_sync_prdy;
wire mul_sync_pvld;
NV_NVDLA_SDP_HLS_sync2data #(.DATA1_WIDTH(16 ),.DATA2_WIDTH(33 )) x_mul_sync2data (
   .chn1_en (!cfg_mul_bypass & cfg_mul_src) //|< ?
  ,.chn2_en (!cfg_mul_bypass) //|< i
  ,.chn1_in_pvld (mul_op_pvld) //|< i
  ,.chn1_in_prdy (mul_op_prdy) //|> o
  ,.chn2_in_pvld (alu_out_pvld) //|< i
  ,.chn2_in_prdy (alu_out_srdy) //|> w
  ,.chn_out_pvld (mul_sync_pvld) //|> w
  ,.chn_out_prdy (mul_sync_prdy) //|< w
  ,.data1_in (chn_mul_op[15:0]) //|< i
  ,.data2_in (alu_data_out[32:0]) //|< i
  ,.data1_out (mul_op_sync[15:0]) //|> w
  ,.data2_out (mul_data_sync[32:0]) //|> w
  );
assign bypass_trt = cfg_mul_prelu & !mul_data_sync[33 -1];
assign mul_op_in[15:0] = (cfg_mul_src == 0 ) ? cfg_mul_op[15:0] : mul_op_sync[15:0];
assign mul_data_in[32:0] = mul_data_sync[32:0];
NV_NVDLA_SDP_HLS_prelu #(.IN_WIDTH(33 ),.OUT_WIDTH(49 ),.OP_WIDTH(16 )) x_mul_prelu (
   .cfg_prelu_en (cfg_mul_prelu) //|< i
  ,.data_in (mul_data_in[32:0]) //|< w
  ,.op_in (mul_op_in[15:0]) //|< w
  ,.data_out (mul_prelu_out[48:0]) //|> w
  );
NV_NVDLA_SDP_HLS_X_INT_MUL_pipe_p1 pipe_p1 (
   .nvdla_core_clk (nvdla_core_clk) //|< i
  ,.nvdla_core_rstn (nvdla_core_rstn) //|< i
  ,.bypass_trt (bypass_trt) //|< w
  ,.mul_final_prdy (mul_final_prdy) //|< w
  ,.mul_prelu_out (mul_prelu_out[48:0]) //|< w
  ,.mul_sync_pvld (mul_sync_pvld) //|< w
  ,.bypass_trt_reg (bypass_trt_reg) //|> w
  ,.mul_data_final (mul_data_final[48:0]) //|> w
  ,.mul_final_pvld (mul_final_pvld) //|> w
  ,.mul_sync_prdy (mul_sync_prdy) //|> w
  );
assign alu_out_prdy = cfg_mul_bypass ? mul_out_prdy : alu_out_srdy;
assign mul_final_prdy = cfg_mul_bypass ? 1'b1 : mul_out_prdy;
assign mul_out_pvld = cfg_mul_bypass ? alu_out_pvld : mul_final_pvld;
assign bypass_trt_out = cfg_mul_bypass ? 1'b0 : bypass_trt_reg;
assign mul_data_out[48:0] = cfg_mul_bypass ? {{16{alu_data_out[32]}}, alu_data_out[32:0]} : mul_data_final[48:0];
endmodule // NV_NVDLA_SDP_HLS_X_int_mul
// **************************************************************************************************************
// Generated by ::pipe -m -bc -rand none -is {mul_data_final[48:0],bypass_trt_reg} (mul_final_pvld,mul_final_prdy) <= {mul_prelu_out[48:0],bypass_trt} (mul_sync_pvld,mul_sync_prdy)
// **************************************************************************************************************
module NV_NVDLA_SDP_HLS_X_INT_MUL_pipe_p1 (
   nvdla_core_clk
  ,nvdla_core_rstn
  ,bypass_trt
  ,mul_final_prdy
  ,mul_prelu_out
  ,mul_sync_pvld
  ,bypass_trt_reg
  ,mul_data_final
  ,mul_final_pvld
  ,mul_sync_prdy
  );
input nvdla_core_clk;
input nvdla_core_rstn;
input bypass_trt;
input mul_final_prdy;
input [48:0] mul_prelu_out;
input mul_sync_pvld;
output bypass_trt_reg;
output [48:0] mul_data_final;
output mul_final_pvld;
output mul_sync_prdy;
reg bypass_trt_reg;
reg [48:0] mul_data_final;
reg mul_final_pvld;
reg mul_sync_prdy;
reg [49:0] p1_pipe_data;
reg p1_pipe_ready;
reg p1_pipe_ready_bc;
reg p1_pipe_valid;
reg p1_skid_catch;
reg [49:0] p1_skid_data;
reg [49:0] p1_skid_pipe_data;
reg p1_skid_pipe_ready;
reg p1_skid_pipe_valid;
reg p1_skid_ready;
reg p1_skid_ready_flop;
reg p1_skid_valid;
//## pipe (1) skid buffer
always @(
  mul_sync_pvld
  or p1_skid_ready_flop
  or p1_skid_pipe_ready
  or p1_skid_valid
  ) begin
  p1_skid_catch = mul_sync_pvld && p1_skid_ready_flop && !p1_skid_pipe_ready;
  p1_skid_ready = (p1_skid_valid)? p1_skid_pipe_ready : !p1_skid_catch;
end
always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
  if (!nvdla_core_rstn) begin
    p1_skid_valid <= 1'b0;
    p1_skid_ready_flop <= 1'b1;
    mul_sync_prdy <= 1'b1;
  end else begin
  p1_skid_valid <= (p1_skid_valid)? !p1_skid_pipe_ready : p1_skid_catch;
  p1_skid_ready_flop <= p1_skid_ready;
  mul_sync_prdy <= p1_skid_ready;
  end
end
always @(posedge nvdla_core_clk) begin
// VCS sop_coverage_off start
  p1_skid_data <= (p1_skid_catch)? {mul_prelu_out[48:0],bypass_trt} : p1_skid_data;
// VCS sop_coverage_off end
end
always @(
  p1_skid_ready_flop
  or mul_sync_pvld
  or p1_skid_valid
  or mul_prelu_out
  or bypass_trt
  or p1_skid_data
  ) begin
  p1_skid_pipe_valid = (p1_skid_ready_flop)? mul_sync_pvld : p1_skid_valid;
// VCS sop_coverage_off start
  p1_skid_pipe_data = (p1_skid_ready_flop)? {mul_prelu_out[48:0],bypass_trt} : p1_skid_data;
// VCS sop_coverage_off end
end
//## pipe (1) valid-ready-bubble-collapse
always @(
  p1_pipe_ready
  or p1_pipe_valid
  ) begin
  p1_pipe_ready_bc = p1_pipe_ready || !p1_pipe_valid;
end
always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
  if (!nvdla_core_rstn) begin
    p1_pipe_valid <= 1'b0;
  end else begin
  p1_pipe_valid <= (p1_pipe_ready_bc)? p1_skid_pipe_valid : 1'd1;
  end
end
always @(posedge nvdla_core_clk) begin
// VCS sop_coverage_off start
  p1_pipe_data <= (p1_pipe_ready_bc && p1_skid_pipe_valid)? p1_skid_pipe_data : p1_pipe_data;
// VCS sop_coverage_off end
end
always @(
  p1_pipe_ready_bc
  ) begin
  p1_skid_pipe_ready = p1_pipe_ready_bc;
end
//## pipe (1) output
always @(
  p1_pipe_valid
  or mul_final_prdy
  or p1_pipe_data
  ) begin
  mul_final_pvld = p1_pipe_valid;
  p1_pipe_ready = mul_final_prdy;
  {mul_data_final[48:0],bypass_trt_reg} = p1_pipe_data;
end
//## pipe (1) assertions/testpoints
`ifndef VIVA_PLUGIN_PIPE_DISABLE_ASSERTIONS
wire p1_assert_clk = nvdla_core_clk;
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML
// spyglass disable_block STARC-2.10.3.2a
// spyglass disable_block STARC05-2.1.3.1
// spyglass disable_block STARC-2.1.4.6
// spyglass disable_block W116
// spyglass disable_block W154
// spyglass disable_block W239
// spyglass disable_block W362
// spyglass disable_block WRN_58
// spyglass disable_block WRN_61
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
// VCS coverage off
  nv_assert_no_x #(0,1,0,"No X's allowed on control signals") zzz_assert_no_x_1x (nvdla_core_clk, `ASSERT_RESET, nvdla_core_rstn, (mul_final_pvld^mul_final_prdy^mul_sync_pvld^mul_sync_prdy)); // spyglass disable W504 SelfDeterminedExpr-ML 
// VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML
// spyglass enable_block STARC-2.10.3.2a
// spyglass enable_block STARC05-2.1.3.1
// spyglass enable_block STARC-2.1.4.6
// spyglass enable_block W116
// spyglass enable_block W154
// spyglass enable_block W239
// spyglass enable_block W362
// spyglass enable_block WRN_58
// spyglass enable_block WRN_61
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML
// spyglass disable_block STARC-2.10.3.2a
// spyglass disable_block STARC05-2.1.3.1
// spyglass disable_block STARC-2.1.4.6
// spyglass disable_block W116
// spyglass disable_block W154
// spyglass disable_block W239
// spyglass disable_block W362
// spyglass disable_block WRN_58
// spyglass disable_block WRN_61
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
// VCS coverage off
  nv_assert_hold_throughout_event_interval #(0,1,0,"valid removed before ready") zzz_assert_hold_throughout_event_interval_2x (nvdla_core_clk, `ASSERT_RESET, (mul_sync_pvld && !mul_sync_prdy), (mul_sync_pvld), (mul_sync_prdy)); // spyglass disable W504 SelfDeterminedExpr-ML 
// VCS coverage on
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML
// spyglass enable_block STARC-2.10.3.2a
// spyglass enable_block STARC05-2.1.3.1
// spyglass enable_block STARC-2.1.4.6
// spyglass enable_block W116
// spyglass enable_block W154
// spyglass enable_block W239
// spyglass enable_block W362
// spyglass enable_block WRN_58
// spyglass enable_block WRN_61
`endif // SPYGLASS_ASSERT_ON
`endif
endmodule // NV_NVDLA_SDP_HLS_X_INT_MUL_pipe_p1
